module engine_null_testbench();

	initial begin
		$display("HI!");
	end

endmodule